library verilog;
use verilog.vl_types.all;
entity EDA3_testbench is
end EDA3_testbench;
