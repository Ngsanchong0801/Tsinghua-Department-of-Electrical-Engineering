library verilog;
use verilog.vl_types.all;
entity EDA3_coincharger_vlg_vec_tst is
end EDA3_coincharger_vlg_vec_tst;
